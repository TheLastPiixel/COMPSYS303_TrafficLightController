
module unsaved (
	clk_clk,
	reset_reset_n,
	sdram_pll_clk_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		sdram_pll_clk_clk;
endmodule
